`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module OR(input [15:0] X, input [15:0] Y, output [15:0] Z);
	assign Z = X | Y;
endmodule
