`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module two_comp(input [15:0] X, output [15:0] Y);
	assign Y = ~X+1;

endmodule
