`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module Full_Adder( A, B, Cin, Sum, Cout);
	input  A, B, Cin;
	output Sum, Cout;	
	wire w;
	
	assign w = A ^ B;
	assign Sum = w ^ Cin;
	assign Cout = (A & B) | (w & Cin); 
	
endmodule
