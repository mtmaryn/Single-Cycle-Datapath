`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module sign_extender( input [7:0] in, output wire[15:0] out);
	
	assign out = {{8{in[7]}}, in[7:0]};

endmodule
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////