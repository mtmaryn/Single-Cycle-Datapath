`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module reg_file( A, B, C, Aaddr, Baddr, Caddr, load, clear, clk );
	input  load, clk, clear;
	input  [15:0] C;
	input  [3:0] Aaddr, Baddr, Caddr;
	output [15:0] A, B;
	


endmodule
